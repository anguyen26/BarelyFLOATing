module random25 (output logic [63:0][15:0] MEM);

	assign MEM[0] = 16'b0001111_111_001_100;
	assign MEM[1] = 16'b0100000001_111_010;
	assign MEM[2] = 16'b0001101_001_100_110;
	assign MEM[3] = 16'b0100000010_011_111;
	assign MEM[4] = 16'b010001100_1011_011;
	assign MEM[5] = 16'b01100_11000_110_111;
	assign MEM[6] = 16'b0100001111_000_010;
	assign MEM[7] = 16'b11100_00000100010;
	assign MEM[8] = 16'b1011_1111_0000_0000;
	assign MEM[9] = 16'b0100001111_011_000;
	assign MEM[10] = 16'b01101_00100_101_100;
	assign MEM[11] = 16'b0001100_111_110_100;
	assign MEM[12] = 16'b010001100_1011_100;
	assign MEM[13] = 16'b01101_00000_101_101;
	assign MEM[14] = 16'b0001110_110_111_001;
	assign MEM[15] = 16'b101100001_0011000;
	assign MEM[16] = 16'b101100001_0001000;
	assign MEM[17] = 16'b0001100_010_001_000;
	assign MEM[18] = 16'b0100000011_001_111;
	assign MEM[19] = 16'b101100001_1100100;
	assign MEM[20] = 16'b0100000100_010_010;
	assign MEM[21] = 16'b101100000_1001000;
	assign MEM[22] = 16'b0001101_000_101_100;
	assign MEM[23] = 16'b0100000000_111_100;
	assign MEM[24] = 16'b0100000011_110_000;
	assign MEM[25] = 16'b0100000111_100_000;
	assign MEM[26] = 16'b01101_00000_000_101;
	assign MEM[27] = 16'b0001111_011_001_111;
	assign MEM[28] = 16'b0001101_100_010_010;
	assign MEM[29] = 16'b0100000010_111_000;
	assign MEM[30] = 16'b0100001111_101_001;
	assign MEM[31] = 16'b01100_10000_010_111;
	assign MEM[32] = 16'b0100000000_011_011;
	assign MEM[33] = 16'b0100001100_101_011;
	assign MEM[34] = 16'b0100001100_111_000;
	assign MEM[35] = 16'b010001100_1010_100;
	assign MEM[36] = 16'b0100000001_010_010;
	assign MEM[37] = 16'b101100001_1000100;
	assign MEM[38] = 16'b0100000100_111_111;
	assign MEM[39] = 16'b0001101_100_000_111;
	assign MEM[40] = 16'b0100001010_110_010;
	assign MEM[41] = 16'b0100000001_000_101;
	assign MEM[42] = 16'b0100000000_001_101;
	assign MEM[43] = 16'b0100000111_010_011;
	assign MEM[44] = 16'b0001101_110_100_110;
	assign MEM[45] = 16'b0100001111_001_001;
	assign MEM[46] = 16'b01101_11100_011_100;
	assign MEM[47] = 16'b00100_010_10101001;
	assign MEM[48] = 16'b0001101_011_000_001;
	assign MEM[49] = 16'b0100000100_111_110;
	assign MEM[50] = 16'b0100001010_000_111;
	assign MEM[51] = 16'b0100000011_101_011;
	assign MEM[52] = 16'b0100001111_010_111;
	assign MEM[53] = 16'b0001111_001_010_011;
	assign MEM[54] = 16'b01100_00000_010_101;
	assign MEM[55] = 16'b0100000100_011_010;
	assign MEM[56] = 16'b0100000011_110_001;
	assign MEM[57] = 16'b0001110_010_000_111;
	assign MEM[58] = 16'b0100000010_100_100;
	assign MEM[59] = 16'b0100001100_001_111;
	assign MEM[60] = 16'b0100001010_101_100;
	assign MEM[61] = 16'b0100001111_000_110;
	assign MEM[62] = 16'b0100000001_011_010;
	assign MEM[63] = 16'b0100000011_111_100;
	assign MEM[64] = 16'b11100_00000000000;

endmodule