module random (output logic [15:0] MEM [63:0]);

	assign MEM[0] = 16'b1110000000000011;
	assign MEM[1] = 16'b0001100001000010;
	assign MEM[2] = 16'b0100011101110000;
	assign MEM[3] = 16'b0010000000000001;
	assign MEM[4] = 16'b0010000100000001;
	assign MEM[5] = 16'b0010001100000000;
	assign MEM[6] = 16'b0010010000000111;
	assign MEM[7] = 16'b0100001010011100;
	assign MEM[8] = 16'b1101100000000110;
	assign MEM[9] = 16'b0100010100111000;
	assign MEM[10] = 16'b0100011000001000;
	assign MEM[11] = 16'b0100011000010001;
	assign MEM[12] = 16'b0001110001011011;
	assign MEM[13] = 16'b1110011111111010;
	assign MEM[14] = 16'b0100011000010011;
	assign MEM[15] = 16'b1011111100000000;
	assign MEM[16] = 16'b1110011111111111;

endmodule