module rotate(
    input logic [15:0] value;
    input logic direction;
    input logic [2:0] distance;

